module range(input [7:0] a, output [3:0] y);

   assign y = a[3:0];

endmodule // range
