module add(input [3:0] a,input[3:0] b, output [5:0] p);

   assign p = a+b;

endmodule
