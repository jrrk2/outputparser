module add(input signed [3:0] a, input signed [3:0] b, output [5:0] p);

   assign p = a+b;

endmodule
