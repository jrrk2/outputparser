module junk;

`define assert(prop)
   
   initial
     `assert(property);

endmodule // junk
