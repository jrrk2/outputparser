module rhs(input a,  output [7:0] z);

   assign z[b] = a;

endmodule // query
